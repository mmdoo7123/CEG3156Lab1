library verilog;
use verilog.vl_types.all;
entity fp_shiftright_norm_vlg_vec_tst is
end fp_shiftright_norm_vlg_vec_tst;
