LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY shiftRegister9 IS
    PORT(
        i_clock, i_resetBar : IN  STD_LOGIC;
        i_load              : IN  STD_LOGIC;
        i_shift             : IN  STD_LOGIC; 
        i_data              : IN  STD_LOGIC_VECTOR(8 downto 0);
        o_q                 : OUT STD_LOGIC_VECTOR(7 downto 0)
    );
END shiftRegister9;

ARCHITECTURE structural OF shiftRegister9 IS
    SIGNAL w_shifted, w_next : STD_LOGIC_VECTOR(8 downto 0);
    SIGNAL w_q               : STD_LOGIC_VECTOR(8 downto 0);
    SIGNAL w_enable          : STD_LOGIC;

    COMPONENT enARdFF_2
        PORT(i_resetBar, i_d, i_enable, i_clock : IN STD_LOGIC; o_q, o_qBar : OUT STD_LOGIC);
    END COMPONENT;

    COMPONENT genericMux2to1
        GENERIC (n : integer := 9);
        PORT(i_A, i_B : IN STD_LOGIC_VECTOR(8 downto 0); i_Sel : IN STD_LOGIC; o_Out : OUT STD_LOGIC_VECTOR(8 downto 0));
    END COMPONENT;

BEGIN
    w_shifted <= '0' & w_q(8 downto 1);

    mux_inst: genericMux2to1
        GENERIC MAP (n => 9)
        PORT MAP (i_A => w_shifted, i_B => i_data, i_Sel => i_load, o_Out => w_next);

    w_enable <= i_load OR i_shift;

    gen_bits: FOR i IN 8 DOWNTO 0 GENERATE
        dff_inst: enARdFF_2
            PORT MAP (
                i_resetBar => i_resetBar,
                i_clock    => i_clock,
                i_enable   => w_enable,
                i_d        => w_next(i),
                o_q        => w_q(i),
                o_qBar     => OPEN
            );
    END GENERATE;

    o_q <= w_q(7 downto 0);
END structural;