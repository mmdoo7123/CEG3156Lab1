library verilog;
use verilog.vl_types.all;
entity toplevelmMULT_vlg_vec_tst is
end toplevelmMULT_vlg_vec_tst;
