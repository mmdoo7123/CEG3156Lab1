library verilog;
use verilog.vl_types.all;
entity fpMultiplier_vlg_vec_tst is
end fpMultiplier_vlg_vec_tst;
