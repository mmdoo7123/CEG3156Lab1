library verilog;
use verilog.vl_types.all;
entity exp_counter7_vlg_vec_tst is
end exp_counter7_vlg_vec_tst;
