library verilog;
use verilog.vl_types.all;
entity eightBitRightShift_vlg_vec_tst is
end eightBitRightShift_vlg_vec_tst;
