library verilog;
use verilog.vl_types.all;
entity exp_counter7 is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        i_load7         : in     vl_logic;
        i_inc1          : in     vl_logic;
        i_data          : in     vl_logic_vector(6 downto 0);
        o_REz           : out    vl_logic_vector(6 downto 0)
    );
end exp_counter7;
