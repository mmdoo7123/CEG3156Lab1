library verilog;
use verilog.vl_types.all;
entity fp_multiplier_array_vlg_vec_tst is
end fp_multiplier_array_vlg_vec_tst;
