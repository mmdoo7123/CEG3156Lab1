library verilog;
use verilog.vl_types.all;
entity ShiftRightReg_vlg_vec_tst is
end ShiftRightReg_vlg_vec_tst;
