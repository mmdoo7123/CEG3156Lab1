library verilog;
use verilog.vl_types.all;
entity exp_counter7_vlg_check_tst is
    port(
        o_REz           : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end exp_counter7_vlg_check_tst;
