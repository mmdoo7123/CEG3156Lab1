library verilog;
use verilog.vl_types.all;
entity ControlPathAdder_vlg_vec_tst is
end ControlPathAdder_vlg_vec_tst;
