library verilog;
use verilog.vl_types.all;
entity ControlPath_vlg_vec_tst is
end ControlPath_vlg_vec_tst;
