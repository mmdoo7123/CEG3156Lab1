library verilog;
use verilog.vl_types.all;
entity overflow_underflow_unit_vlg_vec_tst is
end overflow_underflow_unit_vlg_vec_tst;
