library verilog;
use verilog.vl_types.all;
entity expOverUnderUnit_vlg_vec_tst is
end expOverUnderUnit_vlg_vec_tst;
