LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Entity renamed to reflect 8-bit width for the Lab 1 requirements
ENTITY eightBitComparator IS
    PORT(
        i_Ai, i_Bi            : IN    STD_LOGIC_VECTOR(7 downto 0); -- 8-bit inputs
        o_GT, o_LT, o_EQ      : OUT   STD_LOGIC);
END eightBitComparator;

ARCHITECTURE structural OF eightBitComparator IS
    -- Intermediate signals to carry comparison results between bits
    SIGNAL int_GT, int_LT : STD_LOGIC_VECTOR(7 downto 0);
    SIGNAL gnd : STD_LOGIC;

    -- Component for the 1-bit comparator required by lab specs 
    COMPONENT oneBitComparator
    PORT(
        i_GTPrevious, i_LTPrevious    : IN    STD_LOGIC;
        i_Ai, i_Bi                    : IN    STD_LOGIC;
        o_GT, o_LT                    : OUT   STD_LOGIC);
    END COMPONENT;

BEGIN
    gnd <= '0';

    -- MSB Comparison (Bit 7): No previous bits to compare, so we use gnd
    comp7: oneBitComparator
        PORT MAP (i_GTPrevious => gnd, 
                  i_LTPrevious => gnd,
                  i_Ai => i_Ai(7),
                  i_Bi => i_Bi(7),
                  o_GT => int_GT(7),
                  o_LT => int_LT(7));

    -- Middle Bits (6 down to 1): Chain the results from the bit above
    -- Using a generate statement or manual instantiation for structural clarity
    gen_comp: FOR i IN 6 DOWNTO 0 GENERATE
        comp: oneBitComparator
            PORT MAP (i_GTPrevious => int_GT(i+1), 
                      i_LTPrevious => int_LT(i+1),
                      i_Ai => i_Ai(i),
                      i_Bi => i_Bi(i),
                      o_GT => int_GT(i),
                      o_LT => int_LT(i));
    END GENERATE;

    -- Output Driver: The final result is found at the LSB (Bit 0)
    o_GT <= int_GT(0);
    o_LT <= int_LT(0);
    
    -- If it is neither Greater Than nor Less Than, it must be Equal 
    o_EQ <= int_GT(0) NOR int_LT(0);

END structural;