library verilog;
use verilog.vl_types.all;
entity complementReg_vlg_vec_tst is
end complementReg_vlg_vec_tst;
