library verilog;
use verilog.vl_types.all;
entity fourBitRightShift_vlg_vec_tst is
end fourBitRightShift_vlg_vec_tst;
