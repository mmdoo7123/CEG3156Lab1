library verilog;
use verilog.vl_types.all;
entity ExpAdder_vlg_vec_tst is
end ExpAdder_vlg_vec_tst;
