LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY enASdFF_2 IS 
	PORT(
		i_resetBar	: IN	STD_LOGIC;
		i_d		    : IN	STD_LOGIC;
		i_enable	: IN	STD_LOGIC;
		i_clock		: IN	STD_LOGIC;
		o_q, o_qBar	: OUT	STD_LOGIC);
END enASdFF_2;

ARCHITECTURE rtl OF enASdFF_2 IS
	SIGNAL int_q : STD_LOGIC;
BEGIN
oneBitRegister: PROCESS(i_resetBar, i_clock)
BEGIN
	IF (i_resetBar = '0') THEN
		int_q	<= '1'; -- Forces the state to '1' on reset
	ELSIF (rising_edge(i_clock)) THEN
		IF (i_enable = '1') THEN
			int_q	<=	i_d;
		END IF;
	END IF;
END PROCESS oneBitRegister;
	o_q		<=	int_q;
	o_qBar	<=	not(int_q);
END rtl;